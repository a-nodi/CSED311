`define MEM_TO_EX_FORWARD 2'b01
`define WB_TO_EX_FORWARD 2'b10
`define NO_FORWARD 2'b00

module ForwardingUnit(
    ID_EX_rs1,
    ID_EX_rs2,
    EX_MEM_rd,
    MEM_WB_rd,
    EX_MEM_RegWrite,
    MEM_WB_RegWrite,
    ForwardA,
    ForwardB
);

    input [4:0] ID_EX_rs1;
    input [4:0] ID_EX_rs2;
    input [4:0] EX_MEM_rd;
    input [4:0] MEM_WB_rd;
    input EX_MEM_RegWrite;
    input MEM_WB_RegWrite;
    output reg [1:0] ForwardA;
    output reg [1:0] ForwardB;

    always @(*) begin
        // Forward operation of rs1
        if (ID_EX_rs1 != 0 && ID_EX_rs1 == EX_MEM_rd && EX_MEM_RegWrite) begin // MEM stage
            ForwardA = `MEM_TO_EX_FORWARD;
        end
        else if (ID_EX_rs1 != 0 && ID_EX_rs1 == MEM_WB_rd && MEM_WB_RegWrite) begin // WB state
            ForwardA = `WB_TO_EX_FORWARD;
        end
        else begin
            ForwardA = `NO_FORWARD;
        end

        // Forward operation of rs2
        if (ID_EX_rs2 != 0 && ID_EX_rs2 == EX_MEM_rd && EX_MEM_RegWrite) begin // MEM state
            ForwardB = `MEM_TO_EX_FORWARD;
        end
        else if (ID_EX_rs2 != 0 && ID_EX_rs2 == MEM_WB_rd && MEM_WB_RegWrite) begin // WB state
            ForwardB = `WB_TO_EX_FORWARD;
        end
        else begin
            ForwardB = `NO_FORWARD;
        end

    end

endmodule


