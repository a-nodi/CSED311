`include "opcodes.v"

module Control(
    part_of_inst,
    clk,
    reset,
    
)