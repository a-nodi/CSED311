`include "Constants.v"

module TagTable(
    btb_index,
    corresponding_tag
);
    input [`BTB_INDEX_WIDTH - 1:0] btb_index;
    output reg [`TAG_WIDTH - 1:0] corresponding_tag;




endmodule